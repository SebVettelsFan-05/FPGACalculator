//This is only for 8-bits
//Uses state machine

module double_dabble
(
    input [7:0] i_Binary,
    input clk,

    output [7:0] BCD_rep,
    output o_DV
);





endmodule

